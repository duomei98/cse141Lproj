// Code your design here
`include "reg_file.sv"
`include "PC.sv"
`include "instr_ROM.sv"
`include "dat_mem.sv"
`include "alu.sv"
`include "Control.sv"
`include "top_level.sv"