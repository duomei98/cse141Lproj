`include "alu_tb.sv"
